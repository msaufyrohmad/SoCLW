--********************************************
-- Muhammad Saufy Rohmad
-- EE UiTM Shah Alam
-- System on Chip for Lightweight Cryptography
-- saufy@salam.uitm.edu.my
-- control unit module
--********************************************

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity controlunit is
port
(
	I_clk	:in	std_logic;
	I_reset: in std_logic
);
end controlunit;
	
architecture Behavioral of controlunit is
	
begin
	
end Behavioral;
